--------------------------------------------------------------------------------
--! @file log2_tb.vhd
--! @brief Testbench for 8-bit log base 2 calculator
--! @author Lucas Schneider (lucastrschneider@usp.br)
--! @date 2020/06/17
--------------------------------------------------------------------------------

library ieee;
use ieee.numeric_bit.all;

entity log2_tb is
end log2_tb;